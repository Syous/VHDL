library ieee;
use ieee.std_logic_1164.all;

entity exercise3b is
    port
    (
        A, B, C :   in  std_logic;
        F       :   out std_logic
    );
end entity exercise3b;